--Nicholas Schroeder
-- Testbench for 32-bit ALU

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY ALU_TB IS
END ALU_TB;

ARCHITECTURE TEST_BEHAV OF ALU_TB IS
	COMPONENT ALU
		PORT(
			A		: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
			B		: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
			SHAMT	: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
			ALUOP	: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			OVERFLOW	: OUT STD_LOGIC;
			ZERO		: OUT STD_LOGIC;
			R		: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
		);
	END COMPONENT;

	SIGNAL A			: STD_LOGIC_VECTOR(31 DOWNTO 0) := X"00000000";
	SIGNAL B			: STD_LOGIC_VECTOR(31 DOWNTO 0) := X"00000000";
	SIGNAL SHAMT		: STD_LOGIC_VECTOR(4 DOWNTO 0)  := "00000";
	SIGNAL ALUOP		: STD_LOGIC_VECTOR(3 DOWNTO 0)  := "0000";
	SIGNAL OVERFLOW	: STD_LOGIC;
	SIGNAL ZERO		: STD_LOGIC;
	SIGNAL R			: STD_LOGIC_VECTOR(31 DOWNTO 0);

BEGIN

	ALU_0: ALU PORT MAP(
				A		=> A,
				B		=> B,
				SHAMT	=> SHAMT,	
				ALUOP	=> ALUOP,
				OVERFLOW  => OVERFLOW,
				ZERO		=> ZERO,
				R		=> R);
	PROCESS
	BEGIN

	--TEST CASES PULLED FROM: 
		-- http://people.cs.pitt.edu/~don/coe1502/spring00/Unit1/ALUTest/ALU_TestBench.html

	----LOGIC----

	--TEST AND--
	ALUOP 	<= "0000";
	A		<= "01010101010111110101010101011111";
	B		<= "11111111111111111111111111111111";
	
	WAIT FOR 10 NS;
	ASSERT(R = (A AND B)) REPORT "FAILURE_TEST: AND" SEVERITY FAILURE;

	--TEST OR--
	ALUOP	<= "0001";
	A		<= "01010101010101010101010101010101";
	B		<= "10101010101010101010101010101010";

	WAIT FOR 10 NS;
	ASSERT(R = (A OR B)) REPORT "FAILURE_TEST: OR" SEVERITY FAILURE;

	--TEST XOR--
	ALUOP 	<= "0010";
	A		<= "01010101010101010101010101010101";
	B		<= "11111111111111111111111111111111";
	
	WAIT FOR 10 NS;
	ASSERT(R = (A XOR B)) REPORT "FAILURE_TEST: XOR" SEVERITY FAILURE;

	--TEST NOR--
	ALUOP	<= "0011";
	A		<= "01010101010101010101010101010101";
	B		<= X"00000000";
	WAIT FOR 10 NS;
	ASSERT(R = (A NOR B)) REPORT "FAILURE_TEST: NOR" SEVERITY FAILURE;

	----ARITHMETIC----

	--TEST ADD--
	ALUOP	<= "0100";
	A		<= "01111111111111111111111111111111";
	B		<= "00000000000000000000000000000001";

	WAIT FOR 10 NS;
	ASSERT(R = "10000000000000000000000000000000" AND OVERFLOW = '1' AND ZERO = '0')
	REPORT "FAILURE_TEST: ADD (with overflow)" SEVERITY FAILURE;

	--TEST ADDU--
	ALUOP	<= "0101";

	WAIT FOR 10 NS;
	ASSERT(R = "10000000000000000000000000000000" AND OVERFLOW = '0' AND ZERO = '0')
	REPORT "FAILURE_TEST: ADDU" SEVERITY FAILURE;

	--TEST SUB--
	ALUOP	<= "0110";

	WAIT FOR 10 NS;
	ASSERT(R = "01111111111111111111111111111110" AND OVERFLOW = '0' AND ZERO = '0')
	REPORT "FAILURE_TEST: SUB" SEVERITY FAILURE;	

	--TEST SUBU--
	ALUOP	<= "0110";

	WAIT FOR 10 NS;
	ASSERT(R = "01111111111111111111111111111110" AND OVERFLOW = '0' AND ZERO = '0')
	REPORT "FAILURE_TEST: SUBU" SEVERITY FAILURE;	

	--TEST ADD_2--
	A		<= "10000000000000000000000000000000";
	ALUOP	<= "0100";

	WAIT FOR 10 NS;
	ASSERT(R = "10000000000000000000000000000001" AND OVERFLOW = '0' AND ZERO = '0')
	REPORT "FAILURE_TEST: ADD_2" SEVERITY FAILURE;

	--TEST ADDU_2--
	ALUOP	<= "0101";

	WAIT FOR 10 NS;
	ASSERT(R = "10000000000000000000000000000001" AND OVERFLOW = '0' AND ZERO = '0')
	REPORT "FAILURE_TEST: ADDU_2" SEVERITY FAILURE;

	--TEST SUB_2--
	ALUOP	<= "0110";
	
	WAIT FOR 10 NS;
	ASSERT(R = "01111111111111111111111111111111" AND OVERFLOW = '1' AND ZERO = '0')
	REPORT "FAILURE_TEST: SUB_2" SEVERITY FAILURE;

	--TEST SUBU_2--
	ALUOP	<= "0111";

	WAIT FOR 10 NS;
	ASSERT(R = "01111111111111111111111111111111" AND OVERFLOW = '0' AND ZERO = '0')
	REPORT "FAILURE_TEST: SUBU_2" SEVERITY FAILURE;

	--TEST ADD_ZERO--
	ALUOP	<= "0100";
	A		<= "00000000000000000000000000000001";
	B		<= "11111111111111111111111111111111";

	WAIT FOR 10 NS;
	ASSERT(R = "00000000000000000000000000000000" AND OVERFLOW = '0' AND ZERO = '1')
	REPORT "FAILURE_TEST: ADD_ZERO" SEVERITY FAILURE;	

	----COMPARISON----
	
	--TEST SLT--
	ALUOP	<= "1010";
	A		<= "01111111111111111111111111111111";
	B		<= "00000000000000001111111111111111";

	WAIT FOR 10 NS;
	ASSERT(R = "00000000000000000000000000000000") REPORT "FAILURE_TEST: SLT" SEVERITY FAILURE;

	--TEST SLTU--
	ALUOP	<= "1011";

	WAIT FOR 10 NS;
	ASSERT(R = "00000000000000000000000000000000") REPORT "FAILURE_TEST: SLTU" SEVERITY FAILURE;

	--TEST SLT_2--
	ALUOP 	<= "1010";
	A		<= "00000000000000001111111111111111";
	B		<= "01111111111111111111111111111111";

	WAIT FOR 10 NS;
	ASSERT(R = "00000000000000000000000000000001") REPORT "FAILURE_TEST: SLT_2" SEVERITY FAILURE;

	--TEST SLTU_2--
	ALUOP	<= "1011";

	WAIT FOR 10 NS;
	ASSERT(R = "00000000000000000000000000000001") REPORT "FAILURE_TEST: SLTU_2" SEVERITY FAILURE;

	--TEST SLT_3--
	ALUOP	<= "1010";
	B		<= "11111111111111111111111111111111";

	WAIT FOR 10 NS;
	ASSERT(R = "00000000000000000000000000000000") REPORT "FAILURE_TEST: SLT_3" SEVERITY FAILURE;

	--TEST SLTU_3--
	ALUOP	<= "1011";

	WAIT FOR 10 NS;
	ASSERT(R = "00000000000000000000000000000001") REPORT "FAILURE_TEST: SLTU_3" SEVERITY FAILURE;

	----SHIFTER----
	
	--TEST SLL--
	ALUOP	<= "1100";
	A		<= "11110000000000000000000000001111";
	B		<= "00000000000000000000000000000000";
	SHAMT	<= "01001";

	WAIT FOR 10 NS;
	ASSERT(R = "00000000000000000001111000000000") REPORT "FAILURE_TEST: SLL" SEVERITY FAILURE;

	--TEST SRL--
	ALUOP	<= "1110";

	WAIT FOR 10 NS;
	ASSERT(R = "00000000011110000000000000000000") REPORT "FAILURE_TEST: SRL" SEVERITY FAILURE;

	--TEST SRA--
	ALUOP	<= "1111";

	WAIT FOR 10 NS;
	ASSERT(R = "11111111111110000000000000000000") REPORT "FAILURE_TEST: SRA" SEVERITY FAILURE;



	REPORT "TESTING COMPLETE";
	REPORT "ALL TESTS PASSED";

	WAIT;
	END PROCESS;

END TEST_BEHAV;

