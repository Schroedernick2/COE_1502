--Nicholas Schroeder
-- Mult TB

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY MULT_TB IS
END MULT_TB;

ARCHITECTURE TEST OF MULT_TB IS
	COMPONENT MULTIPLIER_32
		PORT(
			MC		: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
			MP		: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
			RESET	: IN STD_LOGIC;
			START	: IN STD_LOGIC;
			CLOCK	: IN STD_LOGIC;
			PRODUCT	: OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
			DONE		: OUT STD_LOGIC
		);
	END COMPONENT;

	SIGNAL MC		: STD_LOGIC_VECTOR(31 DOWNTO 0) := X"00000000";
	SIGNAL MP		: STD_LOGIC_VECTOR(31 DOWNTO 0) := X"00000000";
	SIGNAL RESET	: STD_LOGIC := '0';
	SIGNAL START	: STD_LOGIC;
	SIGNAL CLOCK	: STD_LOGIC;
	SIGNAL DONE	: STD_LOGIC;
	SIGNAL PRODUCT	: STD_LOGIC_VECTOR(63 DOWNTO 0) := X"0000000000000000";

BEGIN
	MULT_0: MULTIPLIER_32 PORT MAP(MC=>MC,MP=>MP,RESET=>RESET,START=>START,CLOCK=>CLOCK,PRODUCT=>PRODUCT,DONE=>DONE);

	CLOCK_GENERATION: PROCESS
	BEGIN
		CLOCK <= '0';
		WAIT FOR 1 NS;
		CLOCK <= '1';
		WAIT FOR 1 NS;
	END PROCESS CLOCK_GENERATION;

	SIMULATE: PROCESS
	BEGIN
		RESET<='1';
		START<='0';
		WAIT FOR 10 NS;
		RESET<='0';
		MC <= X"00000005";
		MP <= X"00000007";
		START<='1';
		WAIT FOR 20 NS;
		START <= '0';
		WAIT UNTIL DONE='1';

		ASSERT(PRODUCT=X"0000000000000023") REPORT "BIG UH-OH!" SEVERITY FAILURE;

		RESET<='1';
		START<='0';
		WAIT FOR 20 NS;
		RESET<='0';
		MC <= X"0000CDCD";
		MP <= X"01000111";
		START<='1';
		WAIT FOR 20 NS;
		START <= '0';
		WAIT UNTIL DONE='1';

		ASSERT(PRODUCT=X"000000CDCDDB779D") REPORT "BIG UH-OH!" SEVERITY FAILURE;

		RESET<='1';
		START<='0';
		WAIT FOR 20 NS;
		RESET<='0';
		MC <= X"FFFFFFFF";
		MP <= X"00000001";
		START<='1';
		WAIT FOR 20 NS;
		START <= '0';
		WAIT UNTIL DONE='1';

		ASSERT(PRODUCT=X"00000000FFFFFFFF") REPORT "BIG UH-OH!" SEVERITY FAILURE;

		RESET<='1';
		START<='0';
		WAIT FOR 20 NS;
		RESET<='0';
		MC <= X"FFFFFFFF";
		MP <= X"00000000";
		START<='1';
		WAIT FOR 20 NS;
		START <= '0';
		WAIT UNTIL DONE='1';

		ASSERT(PRODUCT=X"0000000000000000") REPORT "BIG UH-OH!" SEVERITY FAILURE;

		WAIT;
	END PROCESS SIMULATE;
END;
