--Nicholas Schroeder
-- Top-Level Unit for 32-bit MIPS CPU

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY TOP_LEVEL IS 
END TOP_LEVEL;

ARCHITECTURE BEHAV OF TOP_LEVEL IS
	SIGNAL CLOCK		: STD_LOGIC;
	SIGNAL RESET		: STD_LOGIC;
	SIGNAL MEM_WAIT 	: STD_LOGIC;
	SIGNAL DATA_OUT		: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL MEM_DATA_OUT	: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL MEM_ADDR		: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL MEM_WRITE	: STD_LOGIC;

	COMPONENT CPU
	PORT(
		RESET			: IN STD_LOGIC;
		CLOCK			: IN STD_LOGIC;
		DATA_MEM_ADDR	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		DATA_MEM_READ	: OUT STD_LOGIC;
		DATA_MEM_WRITE	: OUT STD_LOGIC;
		DATA_MEM_OUT	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		DATA_MEM_WAIT	: IN STD_LOGIC;
		DATA_MEM_IN 	: IN STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
	END COMPONENT;

	COMPONENT COE1502_memory
	PORT(
      Clk      : IN     std_logic;
      MemWrite : IN     std_logic;
      addr     : IN     std_logic_vector (31 DOWNTO 0);
      dataIn   : IN     std_logic_vector (31 DOWNTO 0);
      MemWait  : OUT    std_logic;
      dataOut  : OUT    std_logic_vector (31 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	MEM_0: COE1502_memory
		PORT MAP(
			Clk	=> CLOCK,
			MemWrite => MEM_WRITE,
			addr => MEM_ADDR,
			dataIn => MEM_DATA_OUT,
			MemWait => MEM_WAIT,
			dataOut => DATA_OUT
		);

	CPU_0: CPU
		PORT MAP(
			RESET => RESET,
			CLOCK => CLOCK,
			DATA_MEM_ADDR => MEM_ADDR,
			DATA_MEM_WRITE => MEM_WRITE,
			DATA_MEM_OUT => MEM_DATA_OUT,
			DATA_MEM_WAIT => MEM_WAIT,
			DATA_MEM_IN => DATA_OUT
		);

	CLOCK_GENERATION: PROCESS
	BEGIN
		CLOCK <= '0';
		WAIT FOR 1 NS;
		CLOCK <= '1';
		WAIT FOR 1 NS;
	END PROCESS CLOCK_GENERATION;

	PROCESS
	BEGIN
		RESET <= '1';
		WAIT FOR 10 NS;
		RESET <= '0';
		
		WAIT;
	END PROCESS;

END BEHAV;


























