--Nicholas Schroeder
-- ALU Control for 32-bit MIPS CPU

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY ALU_CONTROL IS
	PORT(
		ALU_OP_IN	: IN STD_LOGIC_VECTOR(3 DOWNTO 0);	--FROM CONTROL
		FUNCT		: IN STD_LOGIC_VECTOR(5 DOWNTO 0);	--INSTR[5-0]
		ALU_OP		: OUT STD_LOGIC_VECTOR(3 DOWNTO 0)	
	);
END ALU_CONTROL;

ARCHITECTURE BEHAV OF ALU_CONTROL IS
BEGIN
	PROCESS(ALU_OP_IN)
	BEGIN

		IF(UNSIGNED(ALU_OP_IN) = 0) THEN
			--R_TYPE CHECK FUNCT--
			IF(UNSIGNED(FUNCT) = 36) THEN
				ALU_OP <= "0000";
			END IF;
			
		ELSE
			--I_TYPE CHECK ALU_OP_IN--
			IF(UNSIGNED(ALU_OP_IN) = 1) THEN
				ALU_OP <= "0100";
			ELSIF(UNSIGNED(ALU_OP_IN) = 2) THEN
				ALU_OP <= "0101";
			ELSIF(UNSIGNED(ALU_OP_IN) = 3) THEN
				ALU_OP <= "1010";
			ELSIF(UNSIGNED(ALU_OP_IN) = 4) THEN
				ALU_OP <= "1011";
			ELSIF(UNSIGNED(ALU_OP_IN) = 5) THEN
				ALU_OP <= "0000";
			ELSIF(UNSIGNED(ALU_OP_IN) = 6) THEN
				ALU_OP <= "0001";
			ELSIF(UNSIGNED(ALU_OP_IN) = 7) THEN
				ALU_OP <= "0010";
			ELSIF(UNSIGNED(ALU_OP_IN) = 8) THEN
				ALU_OP <= "0000"; 	-------LUI HANDLE LATER--------
			END IF;
		END IF;

	END PROCESS;

END BEHAV;
