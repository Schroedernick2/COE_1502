--Nicholas Schroeder
-- 4-bit Ripple Carry Adder

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY ADDER_4 IS
	PORT(
		A		: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		B		: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		CIN		: IN STD_LOGIC;
		COUT 	: OUT STD_LOGIC;
		S		: OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END ADDER_4;

ARCHITECTURE BEHAV OF ADDER_4 IS

	COMPONENT FULL_ADDER
		PORT(
			A		: IN STD_LOGIC;
			B		: IN STD_LOGIC;
			CIN		: IN STD_LOGIC;
			COUT	: OUT STD_LOGIC;
			S		: OUT STD_LOGIC
		);
	END COMPONENT;

	SIGNAL C: STD_LOGIC_VECTOR(3 DOWNTO 0) := "0000";
	SIGNAL SUM: STD_LOGIC_VECTOR(3 DOWNTO 0) := "0000";

BEGIN

	FA0: FULL_ADDER PORT MAP(A=>A(0),B=>B(0),CIN=>CIN,COUT=>C(0),S=>SUM(0)); 
	FA1: FULL_ADDER PORT MAP(A=>A(1),B=>B(1),CIN=>C(0),COUT=>C(1),S=>SUM(1)); 
	FA2: FULL_ADDER PORT MAP(A=>A(2),B=>B(2),CIN=>C(1),COUT=>C(2),S=>SUM(2)); 
	FA3: FULL_ADDER PORT MAP(A=>A(3),B=>B(3),CIN=>C(2),COUT=>C(3),S=>SUM(3)); 

	S 		<= SUM;
	COUT 	<= C(3);

END BEHAV;
