--Nicholas Schroeder
-- test bench for main control unit

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY CONTROL_TB IS
END CONTROL_TB;

ARCHITECTURE BEHAV OF CONTROL_TB IS
	COMPONENT CONTROL
		PORT(
			OP_CODE			: IN STD_LOGIC_VECTOR(5 DOWNTO 0);
			ALU_OP			: OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
			REG_DST			: OUT STD_LOGIC;
			REG_WRITE		: OUT STD_LOGIC;
			ALU_SRC_A		: OUT STD_LOGIC;
			ALU_SRC_B		: OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
			PC_SOURCE		: OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
			PC_WRITE_COND	: OUT STD_LOGIC;
			PC_WRITE		: OUT STD_LOGIC;
			I_OR_D			: OUT STD_LOGIC;
			MEM_READ		: OUT STD_LOGIC;
			MEM_WRITE		: OUT STD_LOGIC;
			MEM_TO_REG		: OUT STD_LOGIC;
			IR_WRITE		: OUT STD_LOGIC;
			CLOCK			: IN STD_LOGIC;
			RESET			: IN STD_LOGIC
		);
	END COMPONENT;

			SIGNAL OP_CODE			: STD_LOGIC_VECTOR(5 DOWNTO 0);
			SIGNAL RESET			: STD_LOGIC;
			SIGNAL CLOCK			: STD_LOGIC;
			SIGNAL ALU_OP			: STD_LOGIC_VECTOR(1 DOWNTO 0);
			SIGNAL REG_DST			: STD_LOGIC;
			SIGNAL REG_WRITE		: STD_LOGIC;
			SIGNAL ALU_SRC_A		: STD_LOGIC;
			SIGNAL ALU_SRC_B		: STD_LOGIC_VECTOR(1 DOWNTO 0);
			SIGNAL PC_SOURCE		: STD_LOGIC_VECTOR(1 DOWNTO 0);
			SIGNAL PC_WRITE_COND	: STD_LOGIC;
			SIGNAL PC_WRITE			: STD_LOGIC;
			SIGNAL I_OR_D			: STD_LOGIC;
			SIGNAL MEM_READ			: STD_LOGIC;
			SIGNAL MEM_WRITE		: STD_LOGIC;
			SIGNAL MEM_TO_REG		: STD_LOGIC;
			SIGNAL IR_WRITE			: STD_LOGIC;

BEGIN
	CONTROL_0: CONTROL PORT MAP(
		OP_CODE => OP_CODE,
		ALU_OP => ALU_OP,
		REG_DST => REG_DST,
		REG_WRITE => REG_WRITE,
		ALU_SRC_A => ALU_SRC_A,
		ALU_SRC_B => ALU_SRC_B,
		PC_SOURCE => PC_SOURCE,
		PC_WRITE_COND => PC_WRITE_COND,
		PC_WRITE => PC_WRITE,
		I_OR_D => I_OR_D,
		MEM_READ => MEM_READ,
		MEM_WRITE => MEM_WRITE,
		MEM_TO_REG => MEM_TO_REG,
		IR_WRITE => IR_WRITE,
		CLOCK => CLOCK,
		RESET => RESET);
		
	PROCESS
	BEGIN
		CLOCK <= '0';
		WAIT FOR 1 NS;
		CLOCK <= '1';
		WAIT FOR 1 NS;
	END PROCESS;

	PROCESS
	BEGIN

		OP_CODE <= "000110";
		--OP_CODE <= "100100";

		WAIT;


	END PROCESS;

END BEHAV;
