--Nicholas Schroeder
-- 32-bit Multiplier

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY MULTIPLIER_32 IS
	PORT(
		MC		: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		MP		: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		RESET	: IN STD_LOGIC;
		START 	: IN STD_LOGIC;
		CLOCK	: IN STD_LOGIC;
		PRODUCT	: OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
		DONE		: OUT STD_LOGIC
	);
END MULTIPLIER_32;

ARCHITECTURE MULTIPLY OF MULTIPLIER_32 IS
	SIGNAL ADD_OUT		: STD_LOGIC_VECTOR(63 DOWNTO 0);
	SIGNAL STOP		: STD_LOGIC:='1';
	SIGNAL SHIFT_MP	: STD_LOGIC:='0';
	SIGNAL SHIFT_MC	: STD_LOGIC:='0';
	SIGNAL PROD_WRITE 	: STD_LOGIC:='0';
	SIGNAL LOAD		: STD_LOGIC:='0';
	SIGNAL COUT		: STD_LOGIC:='0';
	SIGNAL MP_CONTENT	: STD_LOGIC_VECTOR(31 DOWNTO 0) := X"00000000";
	SIGNAL MC_CONTENT	: STD_LOGIC_VECTOR(63 DOWNTO 0) := X"0000000000000000";
	SIGNAL PROD_CONTENT	: STD_LOGIC_VECTOR(63 DOWNTO 0) := X"0000000000000000";

	COMPONENT REG_64B 
		PORT(
			D		: IN STD_LOGIC_VECTOR(63 DOWNTO 0);
			CLOCK	: IN STD_LOGIC;
			ENABLE	: IN STD_LOGIC;
			RESET	: IN STD_LOGIC;
			Q		: OUT STD_LOGIC_VECTOR(63 DOWNTO 0)
		);
	END COMPONENT;

	COMPONENT MP_REG
		PORT(
			MP		: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
			START	: IN STD_LOGIC;
			STOP		: IN STD_LOGIC;
			RESET	: IN STD_LOGIC;
			CLOCK	: IN STD_LOGIC;
			SHIFT	: IN STD_LOGIC;
			CONTENT	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
		); 
	END COMPONENT;

	COMPONENT MC_REG
		PORT(
			MC		: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
			START	: IN STD_LOGIC;
			STOP		: IN STD_LOGIC;
			RESET	: IN STD_LOGIC;
			CLOCK	: IN STD_LOGIC;
			SHIFT	: IN STD_LOGIC;
			CONTENT	: OUT STD_LOGIC_VECTOR(63 DOWNTO 0)
		);
	END COMPONENT;

	COMPONENT ADDER_64
		PORT(
			A		: IN STD_LOGIC_VECTOR(63 DOWNTO 0);
			B		: IN STD_LOGIC_VECTOR(63 DOWNTO 0);
			CIN		: IN STD_LOGIC;
			COUT		: OUT STD_LOGIC;
			S		: OUT STD_LOGIC_VECTOR(63 DOWNTO 0)
		);
	END COMPONENT;

	COMPONENT CONTROL
		PORT(
			MP			: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
			CLOCK		: IN STD_LOGIC;
			START		: IN STD_LOGIC;
			RESET		: IN STD_LOGIC;
			PROD_WRITE	: OUT STD_LOGIC;
			SHIFT_MC		: OUT STD_LOGIC;
			LOAD			: OUT STD_LOGIC;
			SHIFT_MP		: OUT STD_LOGIC;
			STOP			: OUT STD_LOGIC
		);
	END COMPONENT;

BEGIN
	PROD_REG: REG_64B 
		PORT MAP(
			D=>ADD_OUT,
			CLOCK=>CLOCK,
			ENABLE=>PROD_WRITE,
			RESET=>RESET,
			Q=>PROD_CONTENT
		);

	ADDER: ADDER_64 PORT MAP(A=>PROD_CONTENT,B=>MC_CONTENT,CIN=>'0',COUT=>COUT,S=>ADD_OUT);

	MC_REG0: MC_REG PORT MAP(MC=>MC,START=>LOAD,STOP=>STOP,RESET=>RESET,CLOCK=>CLOCK,SHIFT=>SHIFT_MC,CONTENT=>MC_CONTENT);

	MP_REG0: MP_REG PORT MAP(MP=>MP,START=>LOAD,STOP=>STOP,RESET=>RESET,CLOCK=>CLOCK,SHIFT=>SHIFT_MP,CONTENT=>MP_CONTENT);
			
	CTRL: CONTROL PORT MAP(MP=>MP_CONTENT,CLOCK=>CLOCK,PROD_WRITE=>PROD_WRITE,SHIFT_MC=>SHIFT_MC,SHIFT_MP=>SHIFT_MP,START=>START,STOP=>STOP,RESET=>RESET,LOAD=>LOAD);

	PRODUCT <= PROD_CONTENT;
	DONE <= STOP;
END ARCHITECTURE MULTIPLY;
