--Nicholas Schroeder
-- 32-bit Register to store ALU output

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY ALU_OUT_REG IS
	PORT(
		REG_IN		: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		REG_OUT		: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		CLOCK		: IN STD_LOGIC
	);
END ALU_OUT_REG;

ARCHITECTURE BEHAV OF ALU_OUT_REG IS
BEGIN
	PROCESS(CLOCK)
	BEGIN
		IF(RISING_EDGE(CLOCK)) THEN
			REG_OUT <= REG_IN;
		END IF;
	END PROCESS;
END BEHAV;
