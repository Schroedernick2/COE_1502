--Nicholas Schroeder
-- ALU Control for 32-bit MIPS CPU

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY ALU_CONTROL IS
	PORT(
		ALU_OP_IN	: IN STD_LOGIC_VECTOR(3 DOWNTO 0);	--FROM CONTROL
		FUNCT		: IN STD_LOGIC_VECTOR(5 DOWNTO 0);	--INSTR[5-0]
		ALU_OP		: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		SHIFT_SRC : OUT STD_LOGIC;
		SHIFTING : OUT STD_LOGIC;
		CLO     : OUT STD_LOGIC
	);
END ALU_CONTROL;

ARCHITECTURE BEHAV OF ALU_CONTROL IS
BEGIN
	PROCESS(ALU_OP_IN)
	BEGIN
	  CLO <= '0';
	  SHIFTING <= '0';
	  SHIFT_SRC <= '0';

		IF(UNSIGNED(ALU_OP_IN) = 0) THEN
			--R_TYPE CHECK FUNCT--
			IF(UNSIGNED(FUNCT) = 32) THEN
				ALU_OP <= "0100";
			ELSIF(UNSIGNED(FUNCT) = 33) THEN
				ALU_OP <= "0101";
			ELSIF(UNSIGNED(FUNCT) = 34) THEN
				ALU_OP <= "0110";
			ELSIF(UNSIGNED(FUNCT) = 35) THEN
				ALU_OP <= "0111";
			ELSIF(UNSIGNED(FUNCT) = 36) THEN
				ALU_OP <= "0000";
			ELSIF(UNSIGNED(FUNCT) = 37) THEN
				ALU_OP <= "0001";
			ELSIF(UNSIGNED(FUNCT) = 38) THEN
				ALU_OP <= "0010";
			ELSIF(UNSIGNED(FUNCT) = 39) THEN
				ALU_OP <= "0011";
			ELSIF(UNSIGNED(FUNCT) = 42) THEN
				ALU_OP <= "1010";
			ELSIF(UNSIGNED(FUNCT) = 43) THEN
				ALU_OP <= "1011";
			ELSIF(UNSIGNED(FUNCT) = 0) THEN
			  ALU_OP <= "1100";
			  SHIFT_SRC <= '0';
			  SHIFTING <= '1';
			ELSIF(UNSIGNED(FUNCT) = 2) THEN
			  ALU_OP <= "1110";
			  SHIFT_SRC <= '0';
			ELSIF(UNSIGNED(FUNCT) = 3) THEN
			  ALU_OP <= "1111";
			  SHIFT_SRC <= '0';
			  SHIFTING <= '1';
			ELSIF(UNSIGNED(FUNCT) = 4) THEN
			  ALU_OP <= "1100";
			  SHIFT_SRC <= '1';
			  SHIFTING <= '1';
			ELSIF(UNSIGNED(FUNCT) = 6) THEN
			  ALU_OP <= "1110";
			  SHIFT_SRC <= '1';
			  SHIFTING <= '1';
			ELSIF(UNSIGNED(FUNCT) = 7) THEN
			  ALU_OP <= "1111";
			  SHIFT_SRC <= '1';
			  SHIFTING <= '1';
			END IF;
			
		ELSIF(UNSIGNED(ALU_OP_IN) = 15) THEN
		  IF(UNSIGNED(FUNCT) = 33) THEN
		    CLO <= '1';
		  END IF;
			
		ELSE
			--I_TYPE CHECK ALU_OP_IN--
			IF(UNSIGNED(ALU_OP_IN) = 1) THEN
				ALU_OP <= "0100";
			ELSIF(UNSIGNED(ALU_OP_IN) = 2) THEN
				ALU_OP <= "0101";
			ELSIF(UNSIGNED(ALU_OP_IN) = 3) THEN
				ALU_OP <= "1010";
			ELSIF(UNSIGNED(ALU_OP_IN) = 4) THEN
				ALU_OP <= "1011";
			ELSIF(UNSIGNED(ALU_OP_IN) = 5) THEN
				ALU_OP <= "0000";
			ELSIF(UNSIGNED(ALU_OP_IN) = 6) THEN
				ALU_OP <= "0001";
			ELSIF(UNSIGNED(ALU_OP_IN) = 7) THEN
				ALU_OP <= "0010";
			ELSIF(UNSIGNED(ALU_OP_IN) = 8) THEN
				ALU_OP <= "0000"; 	-------LUI HANDLE LATER--------
		  ELSIF(UNSIGNED(ALU_OP_IN) = 9) THEN
		    ALU_OP <= "0110";
			END IF;
		END IF;

	END PROCESS;

END BEHAV;
