--Nicholas Schroeder
-- test bench for CPU

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY CPU_TB IS
END CPU_TB;

ARCHITECTURE BEHAV OF CPU_TB IS
	COMPONENT CPU 
		PORT(
			RESET			: IN STD_LOGIC;
			CLOCK			: IN STD_LOGIC;
			DATA_MEM_ADDR	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DATA_MEM_READ	: OUT STD_LOGIC;
			DATA_MEM_WRITE	: OUT STD_LOGIC;
			DATA_MEM_OUT	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			DATA_MEM_WAIT	: IN STD_LOGIC;
			DATA_MEM_IN 	: IN STD_LOGIC_VECTOR(31 DOWNTO 0)
		);
	END COMPONENT;

	SIGNAL RESET			: STD_LOGIC := '0';
	SIGNAL CLOCK			: STD_LOGIC := '0';
	SIGNAL DATA_MEM_ADDR	: STD_LOGIC_VECTOR(31 DOWNTO 0) := X"00000000";
	SIGNAL DATA_MEM_READ	: STD_LOGIC := '0';
	SIGNAL DATA_MEM_WRITE	: STD_LOGIC := '0';
	SIGNAL DATA_MEM_OUT		: STD_LOGIC_VECTOR(31 DOWNTO 0) := X"00000000";
	SIGNAL DATA_MEM_WAIT	: STD_LOGIC := '0';
	SIGNAL DATA_MEM_IN 		: STD_LOGIC_VECTOR(31 DOWNTO 0) := X"00000000";

BEGIN

	CPU_0: CPU PORT MAP(
		RESET => RESET,
		CLOCK => CLOCK,
		DATA_MEM_ADDR => DATA_MEM_ADDR,
		DATA_MEM_READ => DATA_MEM_READ,
		DATA_MEM_WRITE => DATA_MEM_WRITE,
		DATA_MEM_OUT => DATA_MEM_OUT,
		DATA_MEM_WAIT => DATA_MEM_WAIT,
		DATA_MEM_IN	=> DATA_MEM_IN
	);

	PROCESS
	BEGIN
		CLOCK <= '0';
		WAIT FOR 1 NS;
		CLOCK <= '1';
		WAIT FOR 1 NS;
	END PROCESS;

END BEHAV;
