--Nicholas Schroeder
-- Program Counter for 32-bit MIPS CPU

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY PC IS
	PORT(
		CLOCK	: IN STD_LOGIC;
		RESET	: IN STD_LOGIC;
		PC_IN	: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		ENABLE	: IN STD_LOGIC;
		PC_OUT	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END PC;

ARCHITECTURE BEHAV OF PC IS
BEGIN

	PC_PROC: PROCESS(CLOCK,RESET)
	
	VARIABLE TEMP_PC	: STD_LOGIC_VECTOR(31 DOWNTO 0);

	BEGIN
		IF RESET = '1' THEN
			TEMP_PC := X"00000000";
		ELSIF RISING_EDGE(CLOCK) THEN
			IF ENABLE = '1' THEN
				TEMP_PC := PC_IN;
			END IF;
		END IF;

		PC_OUT <= TEMP_PC;

	END PROCESS;
END BEHAV;			
