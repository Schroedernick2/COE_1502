--Nicholas Schroeder
-- MP Reg

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY MP_REG IS
	PORT(
		MP		: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		START	: IN STD_LOGIC;
		STOP	: IN STD_LOGIC;
		RESET	: IN STD_LOGIC;
		CLOCK	: IN STD_LOGIC;
		SHIFT	: IN STD_LOGIC;
		CONTENT	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END MP_REG;

ARCHITECTURE BEHAV OF MP_REG IS
	COMPONENT REG_32B
		PORT(
			D		: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
			CLOCK	: IN STD_LOGIC;
			ENABLE	: IN STD_LOGIC;
			RESET	: IN STD_LOGIC;
			Q		: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
		);
	END COMPONENT;

	SIGNAL ENABLE			: STD_LOGIC;
	SIGNAL DATA				: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL SHIFTED_CONTENT 	: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL Q				: STD_LOGIC_VECTOR(31 DOWNTO 0);

BEGIN

	REG_32B_0: REG_32B PORT MAP(D=>DATA,CLOCK=>CLOCK,ENABLE=>ENABLE,RESET=>RESET,Q=>Q);

	PROCESS(CLOCK,RESET,STOP,START,SHIFT)
	BEGIN

	ENABLE <= (START OR SHIFT) AND (NOT STOP);

	FOR I IN 0 TO 31 LOOP
		IF(I /= 31) THEN
			SHIFTED_CONTENT(I) <= Q(I+1);
		ELSE
			SHIFTED_CONTENT(I) <= '0';
		END IF;
	END LOOP;

	IF(ENABLE ='1') THEN
		IF(SHIFT='0') THEN
			DATA <= MP;
		ELSIF(SHIFT ='1') THEN
			DATA <= SHIFTED_CONTENT;
		END IF;
	END IF;

	CONTENT <= Q;

	END PROCESS;
END BEHAV;
