--Nicholas Schroeder
-- 64-bit Register

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY REG_64B IS
	PORT(
		D		: IN STD_LOGIC_VECTOR(63 DOWNTO 0);
		CLOCK	: IN STD_LOGIC;
		ENABLE	: IN STD_LOGIC;
		RESET	: IN STD_LOGIC;
		Q		: OUT STD_LOGIC_VECTOR(63 DOWNTO 0)
	);
END REG_64B;

ARCHITECTURE BEHAV OF REG_64B IS
	COMPONENT REG_32B
		PORT(
			D		: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
			CLOCK	: IN STD_LOGIC;
			ENABLE	: IN STD_LOGIC;
			RESET	: IN STD_LOGIC;
			Q		: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
		);
	END COMPONENT;

BEGIN

	REG_32B_0: REG_32B PORT MAP(D(31 DOWNTO 0),CLOCK,ENABLE,RESET,Q(31 DOWNTO 0));
	REG_32B_1: REG_32B PORT MAP(D(63 DOWNTO 32),CLOCK,ENABLE,RESET,Q(63 DOWNTO 32));

END BEHAV;
