LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY ADD_TB IS
END ADD_TB;

ARCHITECTURE BEHAV OF ADD_TB IS
COMPONENT ADDER_64
	PORT(
		A		: IN STD_LOGIC_VECTOR(63 DOWNTO 0);
		B		: IN STD_LOGIC_VECTOR(63 DOWNTO 0);
		CIN		: IN STD_LOGIC;
		COUT		: OUT STD_LOGIC;
		S		: OUT STD_LOGIC_VECTOR(63 DOWNTO 0)
	);
END COMPONENT;

SIGNAL A	: STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL B	: STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL CIN: STD_LOGIC;
SIGNAL COUT: STD_LOGIC;
SIGNAL S	: STD_LOGIC_VECTOR(63 DOWNTO 0);

BEGIN

ADD0: ADDER_64 PORT MAP(A=>A,B=>B,CIN=>CIN,COUT=>COUT,S=>S);
PROCESS
BEGIN
A <= X"000000073E5DE1C7";
B <= X"0000000000000001";
CIN <= '0';

WAIT FOR 10 NS;

ASSERT(S=X"000000073E5DE1C8") REPORT "FUCK" SEVERITY FAILURE;
END PROCESS;
END BEHAV;
