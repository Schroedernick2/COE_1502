--Nicholas Schroeder
-- 4-bit Register

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY REG_4B IS
	PORT(
		D		: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		CLOCK	: IN STD_LOGIC;
		ENABLE	: IN STD_LOGIC;
		RESET	: IN STD_LOGIC;
		Q		: OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END REG_4B;

ARCHITECTURE BEHAV OF REG_4B IS
	COMPONENT REG_1B
		PORT(
			D		: IN STD_LOGIC;
			CLOCK	: IN STD_LOGIC;
			ENABLE	: IN STD_LOGIC;
			RESET	: IN STD_LOGIC;
			Q		: OUT STD_LOGIC
		);
	END COMPONENT;

BEGIN

	REG_1B_0:	REG_1B PORT MAP(D(0),CLOCK,ENABLE,RESET,Q(0));
	REG_1B_1: REG_1B PORT MAP(D(1),CLOCK,ENABLE,RESET,Q(1));
	REG_1B_2:	REG_1B PORT MAP(D(2),CLOCK,ENABLE,RESET,Q(2));
	REG_1B_3: REG_1B PORT MAP(D(3),CLOCK,ENABLE,RESET,Q(3));

END BEHAV;
