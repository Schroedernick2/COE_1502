--Nicholas Schroeder
-- Instruction Register for MIPS 32-bit CPU

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY INSTRUCTION_REG IS
	PORT(
		MEM_DATA		: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		IR_WRITE		: IN STD_LOGIC;
		CLOCK			: IN STD_LOGIC;
		IR_OUT			: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END INSTRUCTION_REG;

ARCHITECTURE BEHAV OF INSTRUCTION_REG IS
BEGIN
	PROCESS(CLOCK,MEM_DATA,IR_WRITE)
	BEGIN
		IF(RISING_EDGE(CLOCK) AND IR_WRITE = '1') THEN
			IR_OUT <= MEM_DATA;
		END IF;
	END PROCESS;
END BEHAV;
