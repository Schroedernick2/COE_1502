LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY REGISTER_FILE_TB IS
END REGISTER_FILE_TB;

ARCHITECTURE BEHAV OF REGISTER_FILE_TB IS

COMPONENT REGISTER_FILE
	PORT(
		CLOCK			: IN STD_LOGIC;
		REG_READ_1_ADDR	: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		REG_READ_2_ADDR	: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		REG_WRITE_ADDR		: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		REG_WRITE			: IN STD_LOGIC;
		REG_WRITE_DATA		: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		REG_READ_1_DATA	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		REG_READ_2_DATA	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

	SIGNAL CLOCK			: STD_LOGIC;
	SIGNAL REG_READ_1_ADDR	: STD_LOGIC_VECTOR(4 DOWNTO 0);
	SIGNAL REG_READ_2_ADDR	: STD_LOGIC_VECTOR(4 DOWNTO 0);
	SIGNAL REG_WRITE_ADDR	: STD_LOGIC_VECTOR(4 DOWNTO 0);
	SIGNAL REG_WRITE		: STD_LOGIC;
	SIGNAL REG_WRITE_DATA	: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL REG_READ_1_DATA	: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL REG_READ_2_DATA	: STD_LOGIC_VECTOR(31 DOWNTO 0);

BEGIN

	RF1: REGISTER_FILE PORT MAP(
		CLOCK=>CLOCK,
		REG_READ_1_ADDR => REG_READ_1_ADDR,
		REG_READ_2_ADDR => REG_READ_2_ADDR,
		REG_WRITE_ADDR => REG_WRITE_ADDR,
		REG_WRITE => REG_WRITE,
		REG_WRITE_DATA => REG_WRITE_DATA,
		REG_READ_1_DATA => REG_READ_1_DATA,
		REG_READ_2_DATA => REG_READ_2_DATA);

	CLOCK_GENERATION: PROCESS
	BEGIN
		CLOCK <= '0';
		WAIT FOR 1 NS;
		CLOCK <= '1';
		WAIT FOR 1 NS;
	END PROCESS CLOCK_GENERATION;

	PROCESS 
	BEGIN
		
	REG_READ_1_ADDR <= "00001";
	REG_READ_2_ADDR <= "00010";

	REG_WRITE_ADDR <= "00001";
	REG_WRITE_DATA <= X"0000FFFF";
	REG_WRITE <= '1';

	WAIT FOR 3 NS;
	REG_WRITE <= '0';	

	WAIT FOR 10 NS;

	REG_WRITE_ADDR <= "00010";
	REG_WRITE_DATA <= X"00000022";
	REG_WRITE <= '1';

	WAIT FOR 2 NS;

	REG_WRITE_ADDR <= "00011";

	WAIT FOR 5 NS;

	REG_WRITE <= '0';

	WAIT FOR 10 NS;

	REG_READ_1_ADDR <= "00011";

	WAIT FOR 10 NS;

	END PROCESS;

END BEHAV;
