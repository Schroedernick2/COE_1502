--Nicholas Schroeder
-- Memory Data Register for MIPS 32-bit CPU

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY MEMORY_REG IS
	PORT(
		MEM_DATA		: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		READ    : IN STD_LOGIC;
		CLOCK			: IN STD_LOGIC;
		MR_OUT			: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END MEMORY_REG;

ARCHITECTURE BEHAV OF MEMORY_REG IS
BEGIN
	PROCESS(CLOCK,MEM_DATA)
	BEGIN
	    IF(READ = '1') THEN
			   MR_OUT <= MEM_DATA;
			END IF;
	END PROCESS;
END BEHAV;
