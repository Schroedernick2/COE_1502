--Nicholas Schroeder
-- Logical Unit for 32-bit ALU

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY LOGICAL_UNIT IS
	PORT(
		A		: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		B		: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		ALUOP	: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		LOGICAL_R : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END LOGICAL_UNIT;

ARCHITECTURE BEHAV OF LOGICAL_UNIT IS
	SIGNAL ANDR	: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL ORR	: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL XORR	: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL NORR	: STD_LOGIC_VECTOR(31 DOWNTO 0);
BEGIN
	ANDR <= A AND B;
	ORR 	<= A OR B;
	XORR <= A XOR B;
	NORR <= A NOR B;

	LOGICAL_R <= 	ANDR WHEN ALUOP = "00" ELSE
				ORR 	WHEN ALUOP = "01" ELSE
				XORR	WHEN ALUOP = "10" ELSE
				NORR;

END BEHAV;
