--Nicholas Schroeder
-- Arithmetic Unit for 32-bit ALU

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY ARITHMETIC_UNIT IS
	PORT(
		ALUOP		: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		A			: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		B			: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		COUT			: OUT STD_LOGIC;
		OVERFLOW		: OUT STD_LOGIC;
		ZERO			: OUT STD_LOGIC;
		ARITHMETIC_R	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END ARITHMETIC_UNIT;

ARCHITECTURE BEHAV OF ARITHMETIC_UNIT IS

	SIGNAL B_TEMP	: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL OFL	: STD_LOGIC;
	SIGNAL S		: STD_LOGIC_VECTOR(31 DOWNTO 0);

	COMPONENT ADDER_32
		PORT(
			A		: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
			B		: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
			CIN		: IN STD_LOGIC;
			COUT 	: OUT STD_LOGIC;
			S		: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
			OFL		: OUT STD_LOGIC
		);
	END COMPONENT;

BEGIN

	B_TEMP 			<= B WHEN ALUOP(1) = '0' ELSE NOT(B);
	OVERFLOW		<= OFL AND NOT(ALUOP(0));
	ARITHMETIC_R	<= S;

	ZERO <= NOT(S(31) OR S(30) OR S(29) OR S(28) OR S(27) OR S(26) OR S(25)
                   OR S(24) OR S(23) OR S(22) OR S(21) OR S(20) OR S(19) OR S(18) OR S(17)               
                   OR S(16) OR S(15) OR S(14) OR S(13) OR S(12) OR S(11) OR S(10) OR S(9)                
                   OR S(8) OR S(7) OR S(6) OR S(5) OR S(4) OR S(3) OR S(2) OR S(1) OR S(0));

	U_0: ADDER_32
		PORT MAP(
			A		=> A,
			B		=> B_TEMP,
			CIN		=> ALUOP(1),
			COUT	=> COUT,
			OFL  	=> OFL,
			S		=> S
		);

END BEHAV;






























