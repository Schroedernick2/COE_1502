--Nicholas Schroeder
-- 4-bit Ripple Carry Adder

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY ADDER_4 IS
	PORT(
		A	: IN	STD_LOGIC_VECTOR(3 DOWNTO 0);
		B	: IN	STD_LOGIC_VECTOR(3 DOWNTO 0);
		CIN	: IN STD_LOGIC;
		COUT : OUT STD_LOGIC;
		S	: OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END ADDER_4;

ARCHITECTURE BEHAV OF ADDER_4 IS

	COMPONENT FULL_ADDER
		PORT(
			A	: IN	STD_LOGIC;
			B	: IN STD_LOGIC;
			CIN	: IN STD_LOGIC;
			COUT	: OUT STD_LOGIC;
			S	: OUT STD_LOGIC
		);
	END COMPONENT;

	SIGNAL C: STD_LOGIC_VECTOR(2 DOWNTO 0);

BEGIN
	FA0:	FULL_ADDER PORT MAP(A(0),B(0),CIN,C(0),S(0));
	FA1:	FULL_ADDER PORT MAP(A(1),B(1),C(0),C(1),S(1));
	FA2:	FULL_ADDER PORT MAP(A(2),B(2),C(1),C(2),S(2));
	FA3:	FULL_ADDER PORT MAP(A(3),B(3),C(2),COUT,S(3));
END BEHAV;
